library verilog;
use verilog.vl_types.all;
entity execute_stage_bench is
end execute_stage_bench;
