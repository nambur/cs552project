library verilog;
use verilog.vl_types.all;
entity generatela is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        \Out\           : out    vl_logic
    );
end generatela;
