library verilog;
use verilog.vl_types.all;
entity carryla_bench is
end carryla_bench;
